/*
    -- System Reset Module --
    Author  : Toddler. 
    Email   : 23011211185@stu.xidian.edu.cn
    Encoder : UTF-8
*/

module sys_rst_m (
    input                 s_clk     ,
    input                 s_rst     ,

    output reg [9 : 0]    o_rst_cnt 
);




endmodule // sys_rst_m
